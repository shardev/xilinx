`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:46:14 01/04/2019 
// Design Name: 
// Module Name:    Multiplekser 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Multiplekser(
    input [15:0] iD0,
    input [15:0] iD1,
    input [15:0] iD2,
    input [15:0] iD3,
    input [15:0] iD4,
    input [15:0] iD5,
    input [15:0] iD6,
    input [15:0] iD7,
    input [15:0] iD8,
    input [3:0] iSEL,
    output [15:0] oQ
    );


endmodule
